
package Hello;

   module mkTb();
      rule hello;
         $display("Hello World!");
         $finish;
      endrule
   endmodule

endpackage

